//********************ѧУ��ɽ���Ƽ���ѧ*****************************//
//********************רҵ��������Ϣ��ѧ�뼼��***********************//
//********************������������***********************************//
//********************ָ����ʦ����С��*******************************//
//********************��Ŀ��CNN�㷨��FPGA������ʵ��******************//
//********************���ڣ�2019.06.01*******************************//
//********************δ��������ֹת��*****************************//

module FC_Para_Set1(
	clk,
	rst,
	
	filt1,
	filt2,
	filt3,
	filt4,
	filt5,
	filt6,
	filt7,
	filt8,
	filt9,
	filt10,
	filt11,
	filt12,
	filt13,
	filt14,
	filt15,
	filt16,
	
	bias1,
	bias2,
	bias3,
	bias4,
	bias5,
	bias6,
	bias7,
	bias8,
	bias9,
	bias10,
	bias11,
	bias12,
	bias13,
	bias14,
	bias15,
	bias16
);

input clk;
input rst;

//���16�����ݣ��ֱ������������ÿ�δ���һ�����ݵĲ�����ʵ�ָ���
output reg [111:0] filt1;
output reg [111:0] filt2;
output reg [111:0] filt3;
output reg [111:0] filt4;
output reg [111:0] filt5;
output reg [111:0] filt6;
output reg [111:0] filt7;
output reg [111:0] filt8;
output reg [111:0] filt9;
output reg [111:0] filt10;
output reg [111:0] filt11;
output reg [111:0] filt12;
output reg [111:0] filt13;
output reg [111:0] filt14;
output reg [111:0] filt15;
output reg [111:0] filt16;

output reg [15:0] bias1;
output reg [15:0] bias2;
output reg [15:0] bias3;
output reg [15:0] bias4;
output reg [15:0] bias5;
output reg [15:0] bias6;
output reg [15:0] bias7;
output reg [15:0] bias8;
output reg [15:0] bias9;
output reg [15:0] bias10;
output reg [15:0] bias11;
output reg [15:0] bias12;
output reg [15:0] bias13;
output reg [15:0] bias14;
output reg [15:0] bias15;
output reg [15:0] bias16;

//�������ظ���Ϊ7*7*4����Ľ�
reg [111:0] para1 [6:0];
reg [111:0] para2 [6:0];
reg [111:0] para3 [6:0];
reg [111:0] para4 [6:0];
reg [111:0] para5 [6:0];
reg [111:0] para6 [6:0];
reg [111:0] para7 [6:0];
reg [111:0] para8 [6:0];
reg [111:0] para9 [6:0];
reg [111:0] para10 [6:0];
reg [111:0] para11 [6:0];
reg [111:0] para12 [6:0];
reg [111:0] para13 [6:0];
reg [111:0] para14 [6:0];
reg [111:0] para15 [6:0];
reg [111:0] para16 [6:0];

integer count;
integer line;

always @(posedge clk)
begin
	if(rst) begin
		count = 0;
		line = 1;
		bias1 = 16'h36;
		bias2 = 16'h36;
		bias3 = 16'h36;
		bias4 = 16'h36;
		bias5 = 16'h36;
		bias6 = 16'h36;
		bias7 = 16'h36;
		bias8 = 16'h36;
		bias9 = 16'h36;
		bias10 = 16'h36;
		bias11 = 16'h36;
		bias12 = 16'h36;
		bias13 = 16'h36;
		bias14 = 16'h36;
		bias15 = 16'h36;
		bias16 = 16'h36;
		para1[0][15:0] = 16'h44;
		para2[0][15:0] = 16'h42;
		para3[0][15:0] = 16'h43;
		para4[0][15:0] = 16'h43;
		para5[0][15:0] = 16'h44;
		para6[0][15:0] = 16'h43;
		para7[0][15:0] = 16'h43;
		para8[0][15:0] = 16'h44;
		para9[0][15:0] = 16'h43;
		para10[0][15:0] = 16'h42;
		para11[0][15:0] = 16'h42;
		para12[0][15:0] = 16'h44;
		para13[0][15:0] = 16'h44;
		para14[0][15:0] = 16'h44;
		para15[0][15:0] = 16'h44;
		para16[0][15:0] = 16'h42;
		para1[0][31:16] = 16'h44;
		para2[0][31:16] = 16'h44;
		para3[0][31:16] = 16'h42;
		para4[0][31:16] = 16'h43;
		para5[0][31:16] = 16'h42;
		para6[0][31:16] = 16'h43;
		para7[0][31:16] = 16'h43;
		para8[0][31:16] = 16'h43;
		para9[0][31:16] = 16'h43;
		para10[0][31:16] = 16'h42;
		para11[0][31:16] = 16'h42;
		para12[0][31:16] = 16'h44;
		para13[0][31:16] = 16'h44;
		para14[0][31:16] = 16'h43;
		para15[0][31:16] = 16'h43;
		para16[0][31:16] = 16'h44;
		para1[0][47:32] = 16'h42;
		para2[0][47:32] = 16'h44;
		para3[0][47:32] = 16'h44;
		para4[0][47:32] = 16'h42;
		para5[0][47:32] = 16'h43;
		para6[0][47:32] = 16'h44;
		para7[0][47:32] = 16'h42;
		para8[0][47:32] = 16'h42;
		para9[0][47:32] = 16'h43;
		para10[0][47:32] = 16'h44;
		para11[0][47:32] = 16'h44;
		para12[0][47:32] = 16'h43;
		para13[0][47:32] = 16'h43;
		para14[0][47:32] = 16'h43;
		para15[0][47:32] = 16'h44;
		para16[0][47:32] = 16'h43;
		para1[0][63:48] = 16'h42;
		para2[0][63:48] = 16'h44;
		para3[0][63:48] = 16'h42;
		para4[0][63:48] = 16'h43;
		para5[0][63:48] = 16'h42;
		para6[0][63:48] = 16'h44;
		para7[0][63:48] = 16'h43;
		para8[0][63:48] = 16'h42;
		para9[0][63:48] = 16'h44;
		para10[0][63:48] = 16'h42;
		para11[0][63:48] = 16'h42;
		para12[0][63:48] = 16'h43;
		para13[0][63:48] = 16'h43;
		para14[0][63:48] = 16'h42;
		para15[0][63:48] = 16'h42;
		para16[0][63:48] = 16'h43;
		para1[0][79:64] = 16'h43;
		para2[0][79:64] = 16'h43;
		para3[0][79:64] = 16'h43;
		para4[0][79:64] = 16'h43;
		para5[0][79:64] = 16'h42;
		para6[0][79:64] = 16'h43;
		para7[0][79:64] = 16'h42;
		para8[0][79:64] = 16'h43;
		para9[0][79:64] = 16'h42;
		para10[0][79:64] = 16'h44;
		para11[0][79:64] = 16'h44;
		para12[0][79:64] = 16'h42;
		para13[0][79:64] = 16'h44;
		para14[0][79:64] = 16'h42;
		para15[0][79:64] = 16'h44;
		para16[0][79:64] = 16'h43;
		para1[0][95:80] = 16'h44;
		para2[0][95:80] = 16'h44;
		para3[0][95:80] = 16'h44;
		para4[0][95:80] = 16'h44;
		para5[0][95:80] = 16'h44;
		para6[0][95:80] = 16'h43;
		para7[0][95:80] = 16'h44;
		para8[0][95:80] = 16'h44;
		para9[0][95:80] = 16'h44;
		para10[0][95:80] = 16'h42;
		para11[0][95:80] = 16'h43;
		para12[0][95:80] = 16'h42;
		para13[0][95:80] = 16'h42;
		para14[0][95:80] = 16'h42;
		para15[0][95:80] = 16'h42;
		para16[0][95:80] = 16'h44;
		para1[0][111:96] = 16'h42;
		para2[0][111:96] = 16'h42;
		para3[0][111:96] = 16'h44;
		para4[0][111:96] = 16'h44;
		para5[0][111:96] = 16'h44;
		para6[0][111:96] = 16'h44;
		para7[0][111:96] = 16'h43;
		para8[0][111:96] = 16'h44;
		para9[0][111:96] = 16'h43;
		para10[0][111:96] = 16'h44;
		para11[0][111:96] = 16'h43;
		para12[0][111:96] = 16'h44;
		para13[0][111:96] = 16'h42;
		para14[0][111:96] = 16'h43;
		para15[0][111:96] = 16'h43;
		para16[0][111:96] = 16'h44;
		para1[1][15:0] = 16'h44;
		para2[1][15:0] = 16'h44;
		para3[1][15:0] = 16'h43;
		para4[1][15:0] = 16'h43;
		para5[1][15:0] = 16'h44;
		para6[1][15:0] = 16'h43;
		para7[1][15:0] = 16'h42;
		para8[1][15:0] = 16'h42;
		para9[1][15:0] = 16'h43;
		para10[1][15:0] = 16'h44;
		para11[1][15:0] = 16'h44;
		para12[1][15:0] = 16'h44;
		para13[1][15:0] = 16'h43;
		para14[1][15:0] = 16'h42;
		para15[1][15:0] = 16'h43;
		para16[1][15:0] = 16'h44;
		para1[1][31:16] = 16'h43;
		para2[1][31:16] = 16'h44;
		para3[1][31:16] = 16'h42;
		para4[1][31:16] = 16'h42;
		para5[1][31:16] = 16'h42;
		para6[1][31:16] = 16'h42;
		para7[1][31:16] = 16'h44;
		para8[1][31:16] = 16'h42;
		para9[1][31:16] = 16'h43;
		para10[1][31:16] = 16'h43;
		para11[1][31:16] = 16'h42;
		para12[1][31:16] = 16'h44;
		para13[1][31:16] = 16'h44;
		para14[1][31:16] = 16'h44;
		para15[1][31:16] = 16'h44;
		para16[1][31:16] = 16'h42;
		para1[1][47:32] = 16'h44;
		para2[1][47:32] = 16'h42;
		para3[1][47:32] = 16'h42;
		para4[1][47:32] = 16'h43;
		para5[1][47:32] = 16'h44;
		para6[1][47:32] = 16'h43;
		para7[1][47:32] = 16'h43;
		para8[1][47:32] = 16'h42;
		para9[1][47:32] = 16'h44;
		para10[1][47:32] = 16'h42;
		para11[1][47:32] = 16'h44;
		para12[1][47:32] = 16'h42;
		para13[1][47:32] = 16'h42;
		para14[1][47:32] = 16'h44;
		para15[1][47:32] = 16'h42;
		para16[1][47:32] = 16'h43;
		para1[1][63:48] = 16'h44;
		para2[1][63:48] = 16'h43;
		para3[1][63:48] = 16'h44;
		para4[1][63:48] = 16'h44;
		para5[1][63:48] = 16'h43;
		para6[1][63:48] = 16'h42;
		para7[1][63:48] = 16'h42;
		para8[1][63:48] = 16'h43;
		para9[1][63:48] = 16'h44;
		para10[1][63:48] = 16'h42;
		para11[1][63:48] = 16'h43;
		para12[1][63:48] = 16'h43;
		para13[1][63:48] = 16'h43;
		para14[1][63:48] = 16'h44;
		para15[1][63:48] = 16'h44;
		para16[1][63:48] = 16'h42;
		para1[1][79:64] = 16'h42;
		para2[1][79:64] = 16'h43;
		para3[1][79:64] = 16'h43;
		para4[1][79:64] = 16'h44;
		para5[1][79:64] = 16'h43;
		para6[1][79:64] = 16'h43;
		para7[1][79:64] = 16'h44;
		para8[1][79:64] = 16'h42;
		para9[1][79:64] = 16'h44;
		para10[1][79:64] = 16'h42;
		para11[1][79:64] = 16'h43;
		para12[1][79:64] = 16'h44;
		para13[1][79:64] = 16'h42;
		para14[1][79:64] = 16'h42;
		para15[1][79:64] = 16'h42;
		para16[1][79:64] = 16'h44;
		para1[1][95:80] = 16'h42;
		para2[1][95:80] = 16'h44;
		para3[1][95:80] = 16'h42;
		para4[1][95:80] = 16'h43;
		para5[1][95:80] = 16'h42;
		para6[1][95:80] = 16'h44;
		para7[1][95:80] = 16'h43;
		para8[1][95:80] = 16'h44;
		para9[1][95:80] = 16'h44;
		para10[1][95:80] = 16'h43;
		para11[1][95:80] = 16'h42;
		para12[1][95:80] = 16'h42;
		para13[1][95:80] = 16'h44;
		para14[1][95:80] = 16'h43;
		para15[1][95:80] = 16'h44;
		para16[1][95:80] = 16'h43;
		para1[1][111:96] = 16'h44;
		para2[1][111:96] = 16'h42;
		para3[1][111:96] = 16'h42;
		para4[1][111:96] = 16'h44;
		para5[1][111:96] = 16'h42;
		para6[1][111:96] = 16'h44;
		para7[1][111:96] = 16'h43;
		para8[1][111:96] = 16'h42;
		para9[1][111:96] = 16'h42;
		para10[1][111:96] = 16'h42;
		para11[1][111:96] = 16'h42;
		para12[1][111:96] = 16'h44;
		para13[1][111:96] = 16'h44;
		para14[1][111:96] = 16'h42;
		para15[1][111:96] = 16'h44;
		para16[1][111:96] = 16'h44;
		para1[2][15:0] = 16'h42;
		para2[2][15:0] = 16'h44;
		para3[2][15:0] = 16'h42;
		para4[2][15:0] = 16'h44;
		para5[2][15:0] = 16'h42;
		para6[2][15:0] = 16'h42;
		para7[2][15:0] = 16'h43;
		para8[2][15:0] = 16'h43;
		para9[2][15:0] = 16'h43;
		para10[2][15:0] = 16'h43;
		para11[2][15:0] = 16'h43;
		para12[2][15:0] = 16'h43;
		para13[2][15:0] = 16'h43;
		para14[2][15:0] = 16'h42;
		para15[2][15:0] = 16'h44;
		para16[2][15:0] = 16'h42;
		para1[2][31:16] = 16'h44;
		para2[2][31:16] = 16'h43;
		para3[2][31:16] = 16'h43;
		para4[2][31:16] = 16'h44;
		para5[2][31:16] = 16'h44;
		para6[2][31:16] = 16'h43;
		para7[2][31:16] = 16'h44;
		para8[2][31:16] = 16'h42;
		para9[2][31:16] = 16'h42;
		para10[2][31:16] = 16'h43;
		para11[2][31:16] = 16'h43;
		para12[2][31:16] = 16'h42;
		para13[2][31:16] = 16'h44;
		para14[2][31:16] = 16'h42;
		para15[2][31:16] = 16'h42;
		para16[2][31:16] = 16'h42;
		para1[2][47:32] = 16'h43;
		para2[2][47:32] = 16'h43;
		para3[2][47:32] = 16'h42;
		para4[2][47:32] = 16'h42;
		para5[2][47:32] = 16'h42;
		para6[2][47:32] = 16'h42;
		para7[2][47:32] = 16'h44;
		para8[2][47:32] = 16'h42;
		para9[2][47:32] = 16'h43;
		para10[2][47:32] = 16'h44;
		para11[2][47:32] = 16'h43;
		para12[2][47:32] = 16'h43;
		para13[2][47:32] = 16'h44;
		para14[2][47:32] = 16'h44;
		para15[2][47:32] = 16'h44;
		para16[2][47:32] = 16'h42;
		para1[2][63:48] = 16'h43;
		para2[2][63:48] = 16'h44;
		para3[2][63:48] = 16'h42;
		para4[2][63:48] = 16'h42;
		para5[2][63:48] = 16'h42;
		para6[2][63:48] = 16'h43;
		para7[2][63:48] = 16'h44;
		para8[2][63:48] = 16'h44;
		para9[2][63:48] = 16'h42;
		para10[2][63:48] = 16'h43;
		para11[2][63:48] = 16'h42;
		para12[2][63:48] = 16'h44;
		para13[2][63:48] = 16'h42;
		para14[2][63:48] = 16'h42;
		para15[2][63:48] = 16'h43;
		para16[2][63:48] = 16'h43;
		para1[2][79:64] = 16'h43;
		para2[2][79:64] = 16'h44;
		para3[2][79:64] = 16'h43;
		para4[2][79:64] = 16'h44;
		para5[2][79:64] = 16'h43;
		para6[2][79:64] = 16'h43;
		para7[2][79:64] = 16'h44;
		para8[2][79:64] = 16'h42;
		para9[2][79:64] = 16'h43;
		para10[2][79:64] = 16'h42;
		para11[2][79:64] = 16'h44;
		para12[2][79:64] = 16'h43;
		para13[2][79:64] = 16'h43;
		para14[2][79:64] = 16'h42;
		para15[2][79:64] = 16'h44;
		para16[2][79:64] = 16'h44;
		para1[2][95:80] = 16'h43;
		para2[2][95:80] = 16'h42;
		para3[2][95:80] = 16'h44;
		para4[2][95:80] = 16'h42;
		para5[2][95:80] = 16'h43;
		para6[2][95:80] = 16'h42;
		para7[2][95:80] = 16'h43;
		para8[2][95:80] = 16'h44;
		para9[2][95:80] = 16'h43;
		para10[2][95:80] = 16'h42;
		para11[2][95:80] = 16'h43;
		para12[2][95:80] = 16'h43;
		para13[2][95:80] = 16'h42;
		para14[2][95:80] = 16'h43;
		para15[2][95:80] = 16'h42;
		para16[2][95:80] = 16'h42;
		para1[2][111:96] = 16'h44;
		para2[2][111:96] = 16'h42;
		para3[2][111:96] = 16'h42;
		para4[2][111:96] = 16'h44;
		para5[2][111:96] = 16'h42;
		para6[2][111:96] = 16'h42;
		para7[2][111:96] = 16'h42;
		para8[2][111:96] = 16'h42;
		para9[2][111:96] = 16'h44;
		para10[2][111:96] = 16'h42;
		para11[2][111:96] = 16'h44;
		para12[2][111:96] = 16'h43;
		para13[2][111:96] = 16'h44;
		para14[2][111:96] = 16'h43;
		para15[2][111:96] = 16'h42;
		para16[2][111:96] = 16'h44;
		para1[3][15:0] = 16'h42;
		para2[3][15:0] = 16'h44;
		para3[3][15:0] = 16'h42;
		para4[3][15:0] = 16'h43;
		para5[3][15:0] = 16'h44;
		para6[3][15:0] = 16'h42;
		para7[3][15:0] = 16'h44;
		para8[3][15:0] = 16'h43;
		para9[3][15:0] = 16'h43;
		para10[3][15:0] = 16'h42;
		para11[3][15:0] = 16'h42;
		para12[3][15:0] = 16'h42;
		para13[3][15:0] = 16'h43;
		para14[3][15:0] = 16'h43;
		para15[3][15:0] = 16'h44;
		para16[3][15:0] = 16'h44;
		para1[3][31:16] = 16'h43;
		para2[3][31:16] = 16'h44;
		para3[3][31:16] = 16'h44;
		para4[3][31:16] = 16'h44;
		para5[3][31:16] = 16'h44;
		para6[3][31:16] = 16'h42;
		para7[3][31:16] = 16'h42;
		para8[3][31:16] = 16'h43;
		para9[3][31:16] = 16'h44;
		para10[3][31:16] = 16'h42;
		para11[3][31:16] = 16'h43;
		para12[3][31:16] = 16'h44;
		para13[3][31:16] = 16'h42;
		para14[3][31:16] = 16'h42;
		para15[3][31:16] = 16'h43;
		para16[3][31:16] = 16'h44;
		para1[3][47:32] = 16'h43;
		para2[3][47:32] = 16'h43;
		para3[3][47:32] = 16'h43;
		para4[3][47:32] = 16'h43;
		para5[3][47:32] = 16'h43;
		para6[3][47:32] = 16'h43;
		para7[3][47:32] = 16'h42;
		para8[3][47:32] = 16'h42;
		para9[3][47:32] = 16'h42;
		para10[3][47:32] = 16'h44;
		para11[3][47:32] = 16'h44;
		para12[3][47:32] = 16'h43;
		para13[3][47:32] = 16'h43;
		para14[3][47:32] = 16'h42;
		para15[3][47:32] = 16'h42;
		para16[3][47:32] = 16'h44;
		para1[3][63:48] = 16'h42;
		para2[3][63:48] = 16'h43;
		para3[3][63:48] = 16'h44;
		para4[3][63:48] = 16'h44;
		para5[3][63:48] = 16'h44;
		para6[3][63:48] = 16'h42;
		para7[3][63:48] = 16'h43;
		para8[3][63:48] = 16'h42;
		para9[3][63:48] = 16'h43;
		para10[3][63:48] = 16'h44;
		para11[3][63:48] = 16'h44;
		para12[3][63:48] = 16'h43;
		para13[3][63:48] = 16'h43;
		para14[3][63:48] = 16'h43;
		para15[3][63:48] = 16'h42;
		para16[3][63:48] = 16'h42;
		para1[3][79:64] = 16'h44;
		para2[3][79:64] = 16'h42;
		para3[3][79:64] = 16'h43;
		para4[3][79:64] = 16'h42;
		para5[3][79:64] = 16'h44;
		para6[3][79:64] = 16'h43;
		para7[3][79:64] = 16'h43;
		para8[3][79:64] = 16'h43;
		para9[3][79:64] = 16'h43;
		para10[3][79:64] = 16'h43;
		para11[3][79:64] = 16'h44;
		para12[3][79:64] = 16'h42;
		para13[3][79:64] = 16'h43;
		para14[3][79:64] = 16'h42;
		para15[3][79:64] = 16'h42;
		para16[3][79:64] = 16'h42;
		para1[3][95:80] = 16'h44;
		para2[3][95:80] = 16'h42;
		para3[3][95:80] = 16'h43;
		para4[3][95:80] = 16'h43;
		para5[3][95:80] = 16'h43;
		para6[3][95:80] = 16'h44;
		para7[3][95:80] = 16'h42;
		para8[3][95:80] = 16'h44;
		para9[3][95:80] = 16'h44;
		para10[3][95:80] = 16'h43;
		para11[3][95:80] = 16'h44;
		para12[3][95:80] = 16'h43;
		para13[3][95:80] = 16'h44;
		para14[3][95:80] = 16'h44;
		para15[3][95:80] = 16'h43;
		para16[3][95:80] = 16'h42;
		para1[3][111:96] = 16'h44;
		para2[3][111:96] = 16'h42;
		para3[3][111:96] = 16'h43;
		para4[3][111:96] = 16'h44;
		para5[3][111:96] = 16'h44;
		para6[3][111:96] = 16'h43;
		para7[3][111:96] = 16'h44;
		para8[3][111:96] = 16'h43;
		para9[3][111:96] = 16'h43;
		para10[3][111:96] = 16'h43;
		para11[3][111:96] = 16'h43;
		para12[3][111:96] = 16'h42;
		para13[3][111:96] = 16'h43;
		para14[3][111:96] = 16'h42;
		para15[3][111:96] = 16'h43;
		para16[3][111:96] = 16'h44;
		para1[4][15:0] = 16'h42;
		para2[4][15:0] = 16'h44;
		para3[4][15:0] = 16'h42;
		para4[4][15:0] = 16'h44;
		para5[4][15:0] = 16'h44;
		para6[4][15:0] = 16'h42;
		para7[4][15:0] = 16'h43;
		para8[4][15:0] = 16'h44;
		para9[4][15:0] = 16'h43;
		para10[4][15:0] = 16'h44;
		para11[4][15:0] = 16'h44;
		para12[4][15:0] = 16'h44;
		para13[4][15:0] = 16'h42;
		para14[4][15:0] = 16'h42;
		para15[4][15:0] = 16'h43;
		para16[4][15:0] = 16'h42;
		para1[4][31:16] = 16'h42;
		para2[4][31:16] = 16'h44;
		para3[4][31:16] = 16'h44;
		para4[4][31:16] = 16'h43;
		para5[4][31:16] = 16'h43;
		para6[4][31:16] = 16'h43;
		para7[4][31:16] = 16'h42;
		para8[4][31:16] = 16'h44;
		para9[4][31:16] = 16'h44;
		para10[4][31:16] = 16'h43;
		para11[4][31:16] = 16'h43;
		para12[4][31:16] = 16'h42;
		para13[4][31:16] = 16'h42;
		para14[4][31:16] = 16'h43;
		para15[4][31:16] = 16'h44;
		para16[4][31:16] = 16'h44;
		para1[4][47:32] = 16'h42;
		para2[4][47:32] = 16'h44;
		para3[4][47:32] = 16'h43;
		para4[4][47:32] = 16'h42;
		para5[4][47:32] = 16'h43;
		para6[4][47:32] = 16'h42;
		para7[4][47:32] = 16'h43;
		para8[4][47:32] = 16'h43;
		para9[4][47:32] = 16'h43;
		para10[4][47:32] = 16'h43;
		para11[4][47:32] = 16'h42;
		para12[4][47:32] = 16'h44;
		para13[4][47:32] = 16'h42;
		para14[4][47:32] = 16'h42;
		para15[4][47:32] = 16'h44;
		para16[4][47:32] = 16'h44;
		para1[4][63:48] = 16'h44;
		para2[4][63:48] = 16'h42;
		para3[4][63:48] = 16'h44;
		para4[4][63:48] = 16'h42;
		para5[4][63:48] = 16'h43;
		para6[4][63:48] = 16'h42;
		para7[4][63:48] = 16'h42;
		para8[4][63:48] = 16'h43;
		para9[4][63:48] = 16'h42;
		para10[4][63:48] = 16'h44;
		para11[4][63:48] = 16'h43;
		para12[4][63:48] = 16'h43;
		para13[4][63:48] = 16'h42;
		para14[4][63:48] = 16'h42;
		para15[4][63:48] = 16'h44;
		para16[4][63:48] = 16'h44;
		para1[4][79:64] = 16'h43;
		para2[4][79:64] = 16'h42;
		para3[4][79:64] = 16'h42;
		para4[4][79:64] = 16'h42;
		para5[4][79:64] = 16'h42;
		para6[4][79:64] = 16'h42;
		para7[4][79:64] = 16'h43;
		para8[4][79:64] = 16'h42;
		para9[4][79:64] = 16'h42;
		para10[4][79:64] = 16'h43;
		para11[4][79:64] = 16'h44;
		para12[4][79:64] = 16'h44;
		para13[4][79:64] = 16'h44;
		para14[4][79:64] = 16'h42;
		para15[4][79:64] = 16'h43;
		para16[4][79:64] = 16'h42;
		para1[4][95:80] = 16'h42;
		para2[4][95:80] = 16'h43;
		para3[4][95:80] = 16'h44;
		para4[4][95:80] = 16'h42;
		para5[4][95:80] = 16'h42;
		para6[4][95:80] = 16'h43;
		para7[4][95:80] = 16'h42;
		para8[4][95:80] = 16'h44;
		para9[4][95:80] = 16'h44;
		para10[4][95:80] = 16'h44;
		para11[4][95:80] = 16'h43;
		para12[4][95:80] = 16'h43;
		para13[4][95:80] = 16'h44;
		para14[4][95:80] = 16'h42;
		para15[4][95:80] = 16'h42;
		para16[4][95:80] = 16'h44;
		para1[4][111:96] = 16'h43;
		para2[4][111:96] = 16'h42;
		para3[4][111:96] = 16'h44;
		para4[4][111:96] = 16'h44;
		para5[4][111:96] = 16'h42;
		para6[4][111:96] = 16'h43;
		para7[4][111:96] = 16'h43;
		para8[4][111:96] = 16'h42;
		para9[4][111:96] = 16'h42;
		para10[4][111:96] = 16'h43;
		para11[4][111:96] = 16'h42;
		para12[4][111:96] = 16'h43;
		para13[4][111:96] = 16'h43;
		para14[4][111:96] = 16'h44;
		para15[4][111:96] = 16'h43;
		para16[4][111:96] = 16'h44;
		para1[5][15:0] = 16'h42;
		para2[5][15:0] = 16'h43;
		para3[5][15:0] = 16'h42;
		para4[5][15:0] = 16'h44;
		para5[5][15:0] = 16'h42;
		para6[5][15:0] = 16'h44;
		para7[5][15:0] = 16'h44;
		para8[5][15:0] = 16'h42;
		para9[5][15:0] = 16'h43;
		para10[5][15:0] = 16'h42;
		para11[5][15:0] = 16'h44;
		para12[5][15:0] = 16'h43;
		para13[5][15:0] = 16'h42;
		para14[5][15:0] = 16'h43;
		para15[5][15:0] = 16'h42;
		para16[5][15:0] = 16'h44;
		para1[5][31:16] = 16'h44;
		para2[5][31:16] = 16'h43;
		para3[5][31:16] = 16'h42;
		para4[5][31:16] = 16'h43;
		para5[5][31:16] = 16'h43;
		para6[5][31:16] = 16'h42;
		para7[5][31:16] = 16'h44;
		para8[5][31:16] = 16'h44;
		para9[5][31:16] = 16'h43;
		para10[5][31:16] = 16'h44;
		para11[5][31:16] = 16'h44;
		para12[5][31:16] = 16'h42;
		para13[5][31:16] = 16'h42;
		para14[5][31:16] = 16'h44;
		para15[5][31:16] = 16'h42;
		para16[5][31:16] = 16'h43;
		para1[5][47:32] = 16'h42;
		para2[5][47:32] = 16'h42;
		para3[5][47:32] = 16'h44;
		para4[5][47:32] = 16'h44;
		para5[5][47:32] = 16'h42;
		para6[5][47:32] = 16'h43;
		para7[5][47:32] = 16'h42;
		para8[5][47:32] = 16'h43;
		para9[5][47:32] = 16'h42;
		para10[5][47:32] = 16'h44;
		para11[5][47:32] = 16'h43;
		para12[5][47:32] = 16'h44;
		para13[5][47:32] = 16'h44;
		para14[5][47:32] = 16'h42;
		para15[5][47:32] = 16'h43;
		para16[5][47:32] = 16'h43;
		para1[5][63:48] = 16'h43;
		para2[5][63:48] = 16'h43;
		para3[5][63:48] = 16'h43;
		para4[5][63:48] = 16'h43;
		para5[5][63:48] = 16'h42;
		para6[5][63:48] = 16'h44;
		para7[5][63:48] = 16'h44;
		para8[5][63:48] = 16'h44;
		para9[5][63:48] = 16'h43;
		para10[5][63:48] = 16'h42;
		para11[5][63:48] = 16'h44;
		para12[5][63:48] = 16'h44;
		para13[5][63:48] = 16'h44;
		para14[5][63:48] = 16'h43;
		para15[5][63:48] = 16'h43;
		para16[5][63:48] = 16'h43;
		para1[5][79:64] = 16'h44;
		para2[5][79:64] = 16'h43;
		para3[5][79:64] = 16'h42;
		para4[5][79:64] = 16'h42;
		para5[5][79:64] = 16'h44;
		para6[5][79:64] = 16'h42;
		para7[5][79:64] = 16'h42;
		para8[5][79:64] = 16'h44;
		para9[5][79:64] = 16'h44;
		para10[5][79:64] = 16'h43;
		para11[5][79:64] = 16'h44;
		para12[5][79:64] = 16'h43;
		para13[5][79:64] = 16'h42;
		para14[5][79:64] = 16'h44;
		para15[5][79:64] = 16'h44;
		para16[5][79:64] = 16'h43;
		para1[5][95:80] = 16'h43;
		para2[5][95:80] = 16'h43;
		para3[5][95:80] = 16'h43;
		para4[5][95:80] = 16'h44;
		para5[5][95:80] = 16'h42;
		para6[5][95:80] = 16'h42;
		para7[5][95:80] = 16'h44;
		para8[5][95:80] = 16'h44;
		para9[5][95:80] = 16'h43;
		para10[5][95:80] = 16'h42;
		para11[5][95:80] = 16'h44;
		para12[5][95:80] = 16'h43;
		para13[5][95:80] = 16'h43;
		para14[5][95:80] = 16'h42;
		para15[5][95:80] = 16'h44;
		para16[5][95:80] = 16'h43;
		para1[5][111:96] = 16'h44;
		para2[5][111:96] = 16'h42;
		para3[5][111:96] = 16'h44;
		para4[5][111:96] = 16'h44;
		para5[5][111:96] = 16'h42;
		para6[5][111:96] = 16'h43;
		para7[5][111:96] = 16'h42;
		para8[5][111:96] = 16'h43;
		para9[5][111:96] = 16'h43;
		para10[5][111:96] = 16'h44;
		para11[5][111:96] = 16'h44;
		para12[5][111:96] = 16'h42;
		para13[5][111:96] = 16'h43;
		para14[5][111:96] = 16'h43;
		para15[5][111:96] = 16'h44;
		para16[5][111:96] = 16'h44;
		para1[6][15:0] = 16'h43;
		para2[6][15:0] = 16'h43;
		para3[6][15:0] = 16'h44;
		para4[6][15:0] = 16'h43;
		para5[6][15:0] = 16'h43;
		para6[6][15:0] = 16'h42;
		para7[6][15:0] = 16'h43;
		para8[6][15:0] = 16'h43;
		para9[6][15:0] = 16'h44;
		para10[6][15:0] = 16'h44;
		para11[6][15:0] = 16'h43;
		para12[6][15:0] = 16'h42;
		para13[6][15:0] = 16'h42;
		para14[6][15:0] = 16'h43;
		para15[6][15:0] = 16'h43;
		para16[6][15:0] = 16'h42;
		para1[6][31:16] = 16'h43;
		para2[6][31:16] = 16'h43;
		para3[6][31:16] = 16'h43;
		para4[6][31:16] = 16'h42;
		para5[6][31:16] = 16'h44;
		para6[6][31:16] = 16'h43;
		para7[6][31:16] = 16'h42;
		para8[6][31:16] = 16'h43;
		para9[6][31:16] = 16'h43;
		para10[6][31:16] = 16'h43;
		para11[6][31:16] = 16'h43;
		para12[6][31:16] = 16'h42;
		para13[6][31:16] = 16'h43;
		para14[6][31:16] = 16'h44;
		para15[6][31:16] = 16'h43;
		para16[6][31:16] = 16'h42;
		para1[6][47:32] = 16'h42;
		para2[6][47:32] = 16'h44;
		para3[6][47:32] = 16'h44;
		para4[6][47:32] = 16'h42;
		para5[6][47:32] = 16'h43;
		para6[6][47:32] = 16'h42;
		para7[6][47:32] = 16'h43;
		para8[6][47:32] = 16'h43;
		para9[6][47:32] = 16'h44;
		para10[6][47:32] = 16'h43;
		para11[6][47:32] = 16'h43;
		para12[6][47:32] = 16'h44;
		para13[6][47:32] = 16'h43;
		para14[6][47:32] = 16'h42;
		para15[6][47:32] = 16'h44;
		para16[6][47:32] = 16'h42;
		para1[6][63:48] = 16'h43;
		para2[6][63:48] = 16'h42;
		para3[6][63:48] = 16'h44;
		para4[6][63:48] = 16'h44;
		para5[6][63:48] = 16'h44;
		para6[6][63:48] = 16'h42;
		para7[6][63:48] = 16'h42;
		para8[6][63:48] = 16'h42;
		para9[6][63:48] = 16'h44;
		para10[6][63:48] = 16'h43;
		para11[6][63:48] = 16'h43;
		para12[6][63:48] = 16'h44;
		para13[6][63:48] = 16'h42;
		para14[6][63:48] = 16'h42;
		para15[6][63:48] = 16'h44;
		para16[6][63:48] = 16'h44;
		para1[6][79:64] = 16'h42;
		para2[6][79:64] = 16'h44;
		para3[6][79:64] = 16'h42;
		para4[6][79:64] = 16'h44;
		para5[6][79:64] = 16'h42;
		para6[6][79:64] = 16'h42;
		para7[6][79:64] = 16'h43;
		para8[6][79:64] = 16'h43;
		para9[6][79:64] = 16'h44;
		para10[6][79:64] = 16'h44;
		para11[6][79:64] = 16'h44;
		para12[6][79:64] = 16'h42;
		para13[6][79:64] = 16'h44;
		para14[6][79:64] = 16'h44;
		para15[6][79:64] = 16'h42;
		para16[6][79:64] = 16'h43;
		para1[6][95:80] = 16'h42;
		para2[6][95:80] = 16'h43;
		para3[6][95:80] = 16'h44;
		para4[6][95:80] = 16'h43;
		para5[6][95:80] = 16'h43;
		para6[6][95:80] = 16'h43;
		para7[6][95:80] = 16'h44;
		para8[6][95:80] = 16'h44;
		para9[6][95:80] = 16'h44;
		para10[6][95:80] = 16'h44;
		para11[6][95:80] = 16'h42;
		para12[6][95:80] = 16'h43;
		para13[6][95:80] = 16'h44;
		para14[6][95:80] = 16'h43;
		para15[6][95:80] = 16'h43;
		para16[6][95:80] = 16'h42;
		para1[6][111:96] = 16'h43;
		para2[6][111:96] = 16'h43;
		para3[6][111:96] = 16'h44;
		para4[6][111:96] = 16'h42;
		para5[6][111:96] = 16'h43;
		para6[6][111:96] = 16'h43;
		para7[6][111:96] = 16'h42;
		para8[6][111:96] = 16'h44;
		para9[6][111:96] = 16'h42;
		para10[6][111:96] = 16'h44;
		para11[6][111:96] = 16'h43;
		para12[6][111:96] = 16'h44;
		para13[6][111:96] = 16'h42;
		para14[6][111:96] = 16'h44;
		para15[6][111:96] = 16'h42;
		para16[6][111:96] = 16'h44;
	end
	
	else begin
		if(line<=6) begin
			filt1 = para1[0];
			filt2 = para2[0];
			filt3 = para3[0];
			filt4 = para4[0];
			filt5 = para5[0];
			filt6 = para6[0];
			filt7 = para7[0];
			filt8 = para8[0];
			filt9 = para9[0];
			filt10 = para10[0];
			filt11 = para11[0];
			filt12 = para12[0];
			filt13 = para13[0];
			filt14 = para14[0];
			filt15 = para15[0];
			filt16 = para16[0];
		end
		
		else if(line<=10) begin
			filt1 = para1[1];
			filt2 = para2[1];
			filt3 = para3[1];
			filt4 = para4[1];
			filt5 = para5[1];
			filt6 = para6[1];
			filt7 = para7[1];
			filt8 = para8[1];
			filt9 = para9[1];
			filt10 = para10[1];
			filt11 = para11[1];
			filt12 = para12[1];
			filt13 = para13[1];
			filt14 = para14[1];
			filt15 = para15[1];
			filt16 = para16[1];
		end
		
		else if(line<=14) begin
			filt1 = para1[2];
			filt2 = para2[2];
			filt3 = para3[2];
			filt4 = para4[2];
			filt5 = para5[2];
			filt6 = para6[2];
			filt7 = para7[2];
			filt8 = para8[2];
			filt9 = para9[2];
			filt10 = para10[2];
			filt11 = para11[2];
			filt12 = para12[2];
			filt13 = para13[2];
			filt14 = para14[2];
			filt15 = para15[2];
			filt16 = para16[2];
		end
		
		else if(line<=18) begin
			filt1 = para1[3];
			filt2 = para2[3];
			filt3 = para3[3];
			filt4 = para4[3];
			filt5 = para5[3];
			filt6 = para6[3];
			filt7 = para7[3];
			filt8 = para8[3];
			filt9 = para9[3];
			filt10 = para10[3];
			filt11 = para11[3];
			filt12 = para12[3];
			filt13 = para13[3];
			filt14 = para14[3];
			filt15 = para15[3];
			filt16 = para16[3];
		end
		
		else if(line<=22) begin
			filt1 = para1[4];
			filt2 = para2[4];
			filt3 = para3[4];
			filt4 = para4[4];
			filt5 = para5[4];
			filt6 = para6[4];
			filt7 = para7[4];
			filt8 = para8[4];
			filt9 = para9[4];
			filt10 = para10[4];
			filt11 = para11[4];
			filt12 = para12[4];
			filt13 = para13[4];
			filt14 = para14[4];
			filt15 = para15[4];
			filt16 = para16[4];
		end
		
		else if(line<=26) begin
			filt1 = para1[5];
			filt2 = para2[5];
			filt3 = para3[5];
			filt4 = para4[5];
			filt5 = para5[5];
			filt6 = para6[5];
			filt7 = para7[5];
			filt8 = para8[5];
			filt9 = para9[5];
			filt10 = para10[5];
			filt11 = para11[5];
			filt12 = para12[5];
			filt13 = para13[5];
			filt14 = para14[5];
			filt15 = para15[5];
			filt16 = para16[5];
		end
		
		else if(line<=30) begin
			filt1 = para1[6];
			filt2 = para2[6];
			filt3 = para3[6];
			filt4 = para4[6];
			filt5 = para5[6];
			filt6 = para6[6];
			filt7 = para7[6];
			filt8 = para8[6];
			filt9 = para9[6];
			filt10 = para10[6];
			filt11 = para11[6];
			filt12 = para12[6];
			filt13 = para13[6];
			filt14 = para14[6];
			filt15 = para15[6];
			filt16 = para16[6];
		end
		
		count = count + 1;
		if(count>25) begin
			count = 0;
			line = line + 1;
			if(line>30) line = 1;
 		end
	end
end



endmodule