//********************ѧУ��ɽ���Ƽ���ѧ*****************************//
//********************רҵ��������Ϣ��ѧ�뼼��***********************//
//********************������������***********************************//
//********************ָ����ʦ����С��*******************************//
//********************��Ŀ��CNN�㷨��FPGA������ʵ��******************//
//********************���ڣ�2019.06.01*******************************//
//********************δ��������ֹת��*****************************//


module clk1(
	clk,
	rst,

	in_pic,
	pic_data
);

input clk;
input rst;
input [223:0] in_pic; //��ROM��ȡ��һ������
output reg [223:0] pic_data; //���һ�����ݵ���һ�������

integer count; //ʱ��ͬ��ʹ��

always @(posedge clk)
begin
	if(rst) count = 0;
	
	else begin
		if(count==0) begin
			pic_data = in_pic;
			count = 1;
			//$display("pic_data = %h", pic_data);
		end
		
		else begin
			count = count + 1;
			if(count==26) count = 0; //26�����ڴ���һ��ͼƬ
		end
	end
end

endmodule