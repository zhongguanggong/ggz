//********************ѧУ��ɽ���Ƽ���ѧ*****************************//
//********************רҵ��������Ϣ��ѧ�뼼��***********************//
//********************������������***********************************//
//********************ָ����ʦ����С��*******************************//
//********************��Ŀ��CNN�㷨��FPGA������ʵ��******************//
//********************���ڣ�2019.06.01*******************************//
//********************δ��������ֹת��*****************************//

//�����λ�ź�����
module rst_gen(
	clk,
	rst_0, 
	rst
);

input clk;
input rst_0;  //������λ�ź�
output reg rst; //�����λ�ź�

integer count;  //ͬ���ź�

always @(posedge clk)
begin
	if(rst_0) begin
		count = 0;
		rst   = 1;
	end
	
	else begin
		count = count + 1;
		if(count>9) begin
			rst = 0;
			count = 9;
		end
	end
end

endmodule